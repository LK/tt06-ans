/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`define default_netname none
`define SYM_WIDTH 4
`define CNT_WIDTH 4

`include "encoder.v"
`include "loader.v"

module ans_encoder_top (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  // assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  // assign uio_out = 0;
  // assign uio_oe  = 0;

  assign uio_oe = 8'b00001111;
  assign uio_in[7:6] = 2'b00;
  assign uo_out[7:4] = 4'b0000;

  ans ans_block (
    .in(ui_in[3:0]),
    .out(uo_out[3:0]),
    .cmd(uio_in[1:0]),
    .in_vld(uio_in[2]),
    .in_rdy(uio_out[4]),
    .out_vld(uio_out[5]),
    .out_rdy(uio_in[3]),
    .clk(clk),
    .rst_n(rst_n)
  );

endmodule

module ans (
  input wire [`SYM_WIDTH-1:0] in,
  output reg [`SYM_WIDTH-1:0] out,
  input wire [1:0] cmd,

  input wire in_vld,
  output wire in_rdy,

  output wire out_vld,
  input wire out_rdy,

  input wire clk,
  input wire rst_n
);

wire mode_enc = cmd == 2'b01;
wire mode_dec = cmd == 2'b10;
wire mode_load = cmd == 2'b11;

wire [`CNT_WIDTH-1:0] counts[2**`SYM_WIDTH-1:0];

wire loader_in_rdy;

ans_loader loader (
  .in(in),
  .counts(counts),
  .in_vld(in_vld),
  .in_rdy(loader_in_rdy),
  .clk(mode_load ? clk : 1'b0),
  .rst_n(rst_n)
);

wire encoder_in_rdy;
wire encoder_out_vld;

ans_encoder encoder (
  .in(in),
  .out(out),
  .in_vld(in_vld),
  .in_rdy(encoder_in_rdy),
  .out_vld(encoder_out_vld),
  .out_rdy(out_rdy),
  .clk(mode_enc ? clk : 1'b0),
  .rst_n(rst_n)
);

assign in_rdy = mode_load ? loader_in_rdy : mode_enc ? encoder_in_rdy : 1'b0;
assign out_vld = mode_enc ? encoder_out_vld : 1'b0;

endmodule
